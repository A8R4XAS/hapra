LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY function_81 IS
    PORT (
--missing
    );
END function_81;

ARCHITECTURE rtl OF function_81 IS

    component mux81 is 
        PORT (--missing);
    end component mux81;

begin
--missing
end rtl;